2 module and gate ( input logic a , b , output logic y ) ;
3 assign y = a & b ;
4 endmodule
